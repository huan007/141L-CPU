//This file defines the parameters used in the alu
package definitions;

typedef enum logic[7:0] {
  IMME = 8'b10??????,
  BLT = 8'b110?????,
  BNE = 8'b111?????,

  ADD = 8'b00000???,
  ADDC = 8'b00001???,
  SUB = 8'b00010???,
  SUBC = 8'b00011???,
  LSL = 8'b00100???,
  LSLC = 8'b00101???,
  LSR = 8'b00110???,
  LSRC = 8'b00111???,
  ASR = 8'b01000???,
  NEG = 8'b01001???,
  AND = 8'b01010???,
  OR = 8'b01011???,
  CMP = 8'b01110???,
  LW = 8'b01101???,
  SW = 8'b01100???,
  ALW = 8'b0111110?,
  ASW = 8'b0111111?,
  HALT = 8'b01110000
} op_code;

endpackage // defintions
