//Program Counter (Fetch)
module IF (
	input 	Abs_Jump,
			Rel_Jump,

